library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity IR is
	port (
		pc: in std_logic_vector (31 downto 0);
		instruction: out std_logic_vector (31 downto 0)
	);
end IR;

architecture behavior of IR is
	type data_rom is array (0 to 31) of std_logic_vector (31 downto 0);
	constant rom: data_rom := (
		"10001100000001110000000000010000", -- lw $t7, 16($0)
		"10001100000010000000000000010010", -- lw $t8, 18($0)
		"00000000111010000100100000100000", -- add $t9, $t7, $t8
		"10101100000010010000000000010100", -- sw $t9, 20($0)
		"10001100000010000000000000010000", -- lw $t8, 16($0)
		"00010000111010000000000000000010", -- beq $t7, $t8, 2
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00001000000000000000000000011111", -- jump here 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000" -- here
	);
	begin
		instruction <= rom(to_integer(unsigned(pc(31 downto 2))));
end behavior;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity IR is
	port (
		pc: in std_logic_vector (31 downto 0);
		instruction: out std_logic_vector (31 downto 0)
	);
end IR;

architecture behavior of IR is
	type data_rom is array (31 downto 0) of std_logic_vector (31 downto 0);
	constant rom: data_rom := (
		"00000000000000001000000000000000",
		"01111100000010000000011111000000",
		"00000000011111010000000100000000",
		"00000000000000000000000000000000",
		"00010000000001000000000011100000",
		"00000000110000000000000000000000",
		"10000000000000000000000000000000",
		"00000011111110000000000000000000",
		"00000000011111001111100000000000",
		"00011100000001000000000011000000", 
		"01111000000000100000000000011111",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"10001100011110000000000110000000", 
		"10111111100000000000011100000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"11111111111111111111111111111110"
	);
	begin
		instruction <= rom(to_integer(unsigned(pc)));
end behavior;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity IR is
	port (
		pc: in std_logic_vector (31 downto 0);
		instruction: out std_logic_vector (31 downto 0)
	);
end IR;

architecture behavior of IR is
	type data_rom is array (0 to 31) of std_logic_vector (31 downto 0);
	constant rom: data_rom := (
		"00100000000010000000000000000111",
		"00100000000010010000000000000110",
		"00100000000010000000000000001000",
		"00100000000010010000000000001000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000"
	);
	begin
		instruction <= rom(to_integer(unsigned(pc(31 downto 2))));
end behavior;
